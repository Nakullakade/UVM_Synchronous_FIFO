package fifo_pkg;

`include "uvm_macros.svh" 
import uvm_pkg::*;

`include "fifo_seq_item.sv"
`include "op_monitor.sv"
`include "ip_monitor.sv"
`include "ip_driver.sv"
`include "ip_seqr.sv"
`include "op_agent.sv"
`include "ip_agent.sv"
`include "fifo_scoreboard.sv"
`include "fifo_func_coverage.sv"
`include "fifo_vseqr.sv"
`include "fifo_env.sv"
`include "fifo_seq.sv"
`include "fifo_vseq.sv"
`include "fifo_test.sv"
endpackage:fifo_pkg